library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL; 
use ieee.numeric_std.all;

entity top is
	port(
		clk: in std_logic
	); 
end top;

architecture Behavioral of top is

begin


end Behavioral;

