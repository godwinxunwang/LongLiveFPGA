library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL; 

entity CPU is
	port (
		input: in std_logic_vector(31 downto 0); 
		output: out std_logic_vector(31 downto 0)
	); 
end CPU;

architecture Behavioral of CPU is

begin


end Behavioral;

